module decoder (
  input [2:0] instruction,
  input sw8,

  output logic rst_count,
  output logic hold_count,

  output logic alu_control

  
  );

  endmodule
