module program_counter (
  input Clock,
  input nReset,
  input branch,
  input rst,
  output logic pc
  );

  endmodule
