module picoMIPS (
  input clk,
  input [9:0] SW,
  output logic [7:0] LED 
  );
  endmodule
