`define ADD 2'b 00 // 3b' RAM 8'b xxxxxRAM

`define IMM 2'b 01 // 3'b RAM 8'b --VALUE--

`define MULT 2'b 10// 3'b RAM (pointer to ROM) 8'b -KERNAL--

`define RBAN 2'b 11// 3'b RAM (rst)
